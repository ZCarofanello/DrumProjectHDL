Freq2StepsMult_inst : Freq2StepsMult PORT MAP (
		clock	 => clock_sig,
		dataa	 => dataa_sig,
		result	 => result_sig
	);
